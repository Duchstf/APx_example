
library IEEE;
use IEEE.STD_LOGIC_1164.all;

use work.StdRtlPkg.all;
use work.ApxL1TPkg.all;
use work.MgtPkg.all;

package PrjSpecPkg is

  constant QPLL_CNT_C   : integer := 24;
  constant REFCLK_CNT_C : integer := 16;
  constant MGT_CNT_C    : integer := 54;

  constant L1T_IN_STREAM_CNT_C  : integer := 54;
  constant L1T_OUT_STREAM_CNT_C : integer := 54;

  constant FS_TO_LHC_CLK_FACTOR_C : integer := 8;

  constant SECTOR_CNT_C : integer := 6;

  constant RefClk0CfgImpl_C : tRefClkCfgArr(0 to REFCLK_CNT_C-1) := (
    0      => (enabled => true, sector => 0),
    1      => (enabled => true, sector => 0),
    2      => (enabled => true, sector => 1),
--  3      => (enabled => true, sector => 1),
    4      => (enabled => true, sector => 1),
    5      => (enabled => true, sector => 2),
    6      => (enabled => true, sector => 2),
    7      => (enabled => true, sector => 2),
    8      => (enabled => true, sector => 3),
    9      => (enabled => true, sector => 3),
    10     => (enabled => true, sector => 4),
    11     => (enabled => true, sector => 4),
    12     => (enabled => true, sector => 4),
    13     => (enabled => true, sector => 5),
    14     => (enabled => true, sector => 5),
    15     => (enabled => true, sector => 5),
    others => RefClkCfgOff_C
    );

  constant RefClk1CfgImpl_C : tRefClkCfgArr(0 to REFCLK_CNT_C-1) := (
    0      => (enabled => true, sector => 0),
    1      => (enabled => true, sector => 0),
    2      => (enabled => true, sector => 1),
    -- 3      => (enabled => true, sector => 1),
    4      => (enabled => true, sector => 1),
    5      => (enabled => true, sector => 2),
    6      => (enabled => true, sector => 2),
    7      => (enabled => true, sector => 2),
    8      => (enabled => true, sector => 3),
    9      => (enabled => true, sector => 3),
    10     => (enabled => true, sector => 4),
    11     => (enabled => true, sector => 4),
    12     => (enabled => true, sector => 4),
    13     => (enabled => true, sector => 5),
    14     => (enabled => true, sector => 5),
    15     => (enabled => true, sector => 5),
    others => RefClkCfgOff_C
    );

  constant QpllCfgImpl_C : tQpllCfgArr(0 to QPLL_CNT_C-1) := (
    0      => (enabled => true, refclk0 => 0, refclk1 => -1, sector => 0),
    1      => (enabled => true, refclk0 => 0, refclk1 => -1, sector => 0),
    2      => (enabled => true, refclk0 => 1, refclk1 => -1, sector => 0),
    3      => (enabled => true, refclk0 => 2, refclk1 => -1, sector => 1),
    4      => (enabled => true, refclk0 => 2, refclk1 => -1, sector => 1),
    5      => (enabled => true, refclk0 => 4, refclk1 => -1, sector => 1),
    6      => (enabled => true, refclk0 => 4, refclk1 => -1, sector => 1),
    7      => (enabled => true, refclk0 => 5, refclk1 => -1, sector => 2),
    8      => (enabled => true, refclk0 => 5, refclk1 => -1, sector => 2),
    9      => (enabled => true, refclk0 => 6, refclk1 => -1, sector => 2),
    10     => (enabled => true, refclk0 => 7, refclk1 => -1, sector => 2),
    11     => (enabled => true, refclk0 => 7, refclk1 => -1, sector => 2),
    12     => (enabled => true, refclk0 => 8, refclk1 => -1, sector => 3),
    13     => (enabled => true, refclk0 => 9, refclk1 => -1, sector => 3),
    14     => (enabled => true, refclk0 => 10, refclk1 => -1, sector => 4),
    15     => (enabled => true, refclk0 => 10, refclk1 => -1, sector => 4),
    16     => (enabled => true, refclk0 => 11, refclk1 => -1, sector => 4),
    17     => (enabled => true, refclk0 => 12, refclk1 => -1, sector => 4),
    18     => (enabled => true, refclk0 => 12, refclk1 => -1, sector => 4),
    19     => (enabled => true, refclk0 => 13, refclk1 => -1, sector => 5),
    20     => (enabled => true, refclk0 => 13, refclk1 => -1, sector => 5),
    21     => (enabled => true, refclk0 => 14, refclk1 => -1, sector => 5),
    22     => (enabled => true, refclk0 => 15, refclk1 => -1, sector => 5),
    23     => (enabled => true, refclk0 => 15, refclk1 => -1, sector => 5),
    others => QpllCfgOff_C
    );

  constant MgtCfgImpl_C : tMgtCfgArr(0 to MGT_CNT_C-1) := (
    0  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    1  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    2  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    3  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    4  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    5  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    6  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    7  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    8  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    9  => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    10 => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    11 => (kind => gty_sym_25p78125, sector => 0, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    12 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    13 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    14 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    15 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    16 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    17 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    18 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    19 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    20 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    21 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    22 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    23 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    24 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    25 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    26 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    27 => (kind => gty_sym_25p78125, sector => 1, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    28 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    29 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    30 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    31 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    32 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    33 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    34 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    35 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    36 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    37 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    38 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    39 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    40 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    41 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    42 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    43 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    44 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    45 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    46 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    47 => (kind => gty_sym_25p78125, sector => 2, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    48 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    49 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    50 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    51 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    52 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    53 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --54 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --55 => (kind => gty_sym_25p78125, sector => 3, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    --56 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --57 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --58 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --59 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --60 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --61 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --62 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --63 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --64 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --65 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --66 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --67 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --68 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --69 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --70 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --71 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --72 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --73 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --74 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --75 => (kind => gty_sym_25p78125, sector => 4, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    --76 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --77 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --78 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --79 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --80 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --81 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --82 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --83 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --84 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --85 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --86 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --87 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --88 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --89 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --90 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --91 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --92 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --93 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --94 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),
    --95 => (kind => gty_sym_25p78125, sector => 5, rxLineRate => 25871250, rx_enc => enc_64b66b, txLineRate => 25871250, tx_enc => enc_64b66b),

    others => MgtCfgOff_C
    );

  constant apxL1TCfgArrImpl : tApxL1TCfgArr(0 to L1T_IN_STREAM_CNT_C-1) := (
    0  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    1  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    2  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    3  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    4  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    5  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    6  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    7  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    8  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    9  => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    10 => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    11 => (sector => 0, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),

    12 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    13 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    14 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    15 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    16 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    17 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    18 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    19 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    20 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    21 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    22 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    23 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    24 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    25 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    26 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    27 => (sector => 1, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),

    28 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    29 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    30 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    31 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    32 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    33 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    34 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    35 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    36 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    37 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    38 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    39 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    40 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    41 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    42 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    43 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    44 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    45 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    46 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    47 => (sector => 2, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),

    48 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    49 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    50 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    51 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    52 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    53 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16)
    --54 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --55 => (sector => 3, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),

    --56 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --57 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --58 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --59 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --60 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --61 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --62 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --63 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --64 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --65 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --66 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --67 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --68 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --69 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --70 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --71 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --72 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --73 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --74 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --75 => (sector => 4, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),

    --76 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --77 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --78 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --79 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --80 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --81 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --82 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --83 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --84 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --85 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --86 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --87 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --88 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --89 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --90 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --91 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --92 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --93 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --94 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16),
    --95 => (sector => 5, linkBufKindRx => buf_72b, frameLengthRx => 48, fifoReadLengthRx => 48, fifoHoldLengthRx => 0, crcLengthRx => 16, linkBufKindTx => buf_72b, frameLengthTx => 48, fifoReadLengthTx => 48, fifoHoldLengthTx => 0, crcLengthTx => 16)
    );

end package PrjSpecPkg;
